module orGate(A,B,X);

    input A,B;
    output X;
    or (X,A,B);
    
endmodule