module tb();

  reg [31:0] A,B;
  reg [2:0] ctrl;
  wire [31:0] Result;
  wire Z,N,C,V;
  
  Flags_ALU dut(
    .A(A), .B(B), .ctrl(ctrl), .Result(Result), .Z(Z), .N(N), .C(C), .V(V)
  );

  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0);
  end

  initial begin
    A <= 32'b00000000000000000000000001000110;
    B <= 32'b00000000000000000000000000110010;
    ctrl <= 3'b000;
    #100;
    
    A <= 32'b00000000000000000001000000111100;
    B <= 32'b00000000000000000001000000111100;
    ctrl <= 3'b001;
    #100;

    A <= 32'b10000000000000000000000000000011;
    B <= 32'b10000000000000000000000000000000;
    ctrl <= 3'b000;
    #100;
      
    A <= 32'b01010101010101010101010101010101;
    B <= 32'b10101010101010101010101010101010;
    ctrl <= 3'b010;
    #100;
    
    A <= 32'b00001110000000000000000000000001;
    B <= 32'b00000000000000110000000000001111;
    ctrl <= 3'b011;
    #100;
  end

endmodule