module notGate(A,B);

    input A;
    output B;
    not (B,A);

endmodule